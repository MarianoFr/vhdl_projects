--------------------------- Sequential Code ---------------------------
-- PROCESSES, FUNCTIONS, and PROCEDURES are the only sections of code that are executed
-- sequentially. However, as a whole, any of these blocks is still concurrent with any
-- other statements placed outside it.
-- Sequential statements are only allowed inside PROCESSES, FUNCTIONS, and PROCEDURES,
-- they are: IF, WAIT,CASE, and LOOP. VARIABLES are also only allowed in sequential code
-- FUNCTIONS and PROCEDURES are very similar to PROCESSES, but are intended for 
-- system-level design, here will only address PROCESSES.
--    PROCESS
-- A PROCESS is a sequential section of VHDL code. It is characterized by the presence 
-- of IF, WAIT, CASE, or LOOP, and by a sensitivity list (except when WAIT is
-- used). A PROCESS must be installed in the main code, and is executed every time a
-- signal in the sensitivity list changes (or the condition related to WAIT is fulfilled). Its
-- syntax is shown below. VARIABLES are optional.
-- [label:] PROCESS (sensitivity list)
--    [VARIABLE name type [range] [:= initial_value;]] -- initial value not synthesizable, only taken into consideration in simulations.
-- BEGIN
--    (sequential code)
-- END PROCESS [label];
-- The use of a label is also optional. Its purpose is to improve code readability.
-- To construct a synchronous circuit, monitoring a signal (clock, for example) is
-- necessary.
-- A D-type flip-flop is the most basic building block in sequential logic circuits
-- -------------------------------------------------
-- LIBRARY ieee;
-- USE ieee.std_logic_1164.all;
-- ENTITY dff IS
--    PORT (d, clk, rst: IN STD_LOGIC;
--       q: OUT STD_LOGIC);
-- END dff;
-- ARCHITECTURE behavior OF dff IS
-- BEGIN
--    PROCESS (clk, rst)
--    BEGIN
--       IF (rst='1') THEN
--          q <= '0';
--       ELSIF (clk'EVENT AND clk='1') THEN -- could be achieved with rising-edge
--          q <= d;
--       END IF;
--    END PROCESS;
-- END behavior;
-- -------------------------------------------------
--   Signals and Variables
-- VHDL has two ways of passing non-static values around: by means of a SIGNAL
-- or by means of a VARIABLE. A SIGNAL can be declared in a PACKAGE,
-- ENTITY or ARCHITECTURE (in its declarative part), while a VARIABLE can
-- only be declared inside a piece of sequential code (in a PROCESS, for example).
--
-- The value of a VARIABLE can never be passed out of the PROCESS directly; if
-- necessary, then it must be assigned to a SIGNAL. On the other hand, the update of a
-- VARIABLE is immediate, that is, we can promptly count on its new value in the
-- next line of code. That is not the case with a SIGNAL (when used in a PROCESS),
-- for its new value is generally only guaranteed to be available after the conclusion of
-- the present run of the PROCESS.
-- Finally, recall from section 4.1 that the assignment operator for a SIGNAL is
--‘‘<=’’ (ex.: sig <¼ 5), while for a VARIABLE it is ‘‘:=’’ (ex.: var :¼ 5).
--
-- *************** IF ***************
-- IF conditions THEN assignments;
-- ELSIF conditions THEN assignments;
-- ...
-- ELSE assignments;
-- END IF;
-- *************** WAIT ****************
-- The WAIT statement is similar to the IF, but it can be used in more than one way.
-- When using the WAIT statement the PROCESS cannot have a sensitivity list.
-- There are 3 syntaxes for the WAIT statement.
-- WAIT UNTIL signal_condition;
-- WAIT ON signal1 [, signal2, ... ];
-- WAIT FOR time;
-- WAIT UNTIL works with a single signal, thus it's more appropiate for writing synchronous 
-- code rather than asynchronous. Because there is no sensitivity list, WAIT UNTIL must 
-- be the first statement in the PROCESS block. This block will execute every time the wait 
-- condition is met.
-------------------------------------------
-- PROCESS -- no sensitivity list
-- BEGIN
--    WAIT UNTIL (clk'EVENT AND clk='1');
--    IF (rst='1') THEN
--       output <= "00000000";
--    ELSIF (clk'EVENT AND clk='1') THEN
--       output <= input;
--    END IF;
-- END PROCESS;
-------------------------------------------
-- WAIT ON accepts multiple signals. In the example below, the PROCESS will
-- continue execution whenever a change in rst or clk occurs.
-------------------------------------------
-- PROCESS
-- BEGIN
--    WAIT ON clk, rst;
--    IF (rst = '1') THEN-- activo en alto
--       output <= "00000000";
--    ELSIF (clk'EVENT AND clk='1') THEN
--       output <= input;
--    END IF;
-- END PROCESS;
-------------------------------------------
-- Finally, WAIT FOR is intended for simulation only (waveform generation for
-- testbenches). Example: WAIT FOR 5ns;
--
-- *************** CASE ****************
-- This is another statement for sequential code. The syntax is below.
-- CASE identifier IS
--    WHEN value => assignments;
--    WHEN value => assignments;
--    ...
-- END CASE;
-- Example:
--    CASE control IS
--       WHEN "00" => x<=a; y<=b;
--       WHEN "01" => x<=b; y<=c;
--       WHEN OTHERS => x<="0000"; y<="ZZZZ";
--    END CASE;
--
-- *************** LOOP ****************
-- Because it's a sequential statement, it can only be used within a PROCESS.
-- FOR/LOOP
-- [label:] FOR identifier IN range LOOP
--    (sequential statements)
-- END LOOP [label];
-- WHILE/LOOP
-- [label:] WHILE condition LOOP
--    (sequential statements)
-- END LOOP [label];
-- 
-- Just like with the GENERATE command, limits must be static.
-- WHILE/LOOP
-- WHILE (i < 10) LOOP
--    WAIT UNTIL clk'EVENT AND clk='1';
--    (other statements)
-- END LOOP;
--
-- We can also use an exit clause, similar to a break in c
-- FOR i IN data'RANGE LOOP
--    CASE data(i) IS
--       WHEN '0' => count:=count+1;
--       WHEN OTHERS => EXIT;
--    END CASE;
-- END LOOP;
--
-- A NEXT satemtent also exists to skip one iteration, similar to continue in c.
--
-- FOR i IN 0 TO 15 LOOP
--    NEXT WHEN i=skip; -- jumps to next iteration
--      (...)
-- END LOOP;
--
-- 